//
//      Project:  Aurora Module Generator version 3.0
//
//         Date:  $Date: 2008/07/21 10:19:46 $
//          Tag:  $Name: i+IP+144966 $
//         File:  $RCSfile: frame_check.ejava,v $
//          Rev:  $Revision: 1.1.2.2 $
//
//      Company:  Xilinx
//
//   Disclaimer:  XILINX IS PROVIDING THIS DESIGN, CODE, OR
//                INFORMATION "AS IS" SOLELY FOR USE IN DEVELOPING
//                PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY
//                PROVIDING THIS DESIGN, CODE, OR INFORMATION AS
//                ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE,
//                APPLICATION OR STANDARD, XILINX IS MAKING NO
//                REPRESENTATION THAT THIS IMPLEMENTATION IS FREE
//                FROM ANY CLAIMS OF INFRINGEMENT, AND YOU ARE
//                RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY
//                REQUIRE FOR YOUR IMPLEMENTATION.  XILINX
//                EXPRESSLY DISCLAIMS ANY WARRANTY WHATSOEVER WITH
//                RESPECT TO THE ADEQUACY OF THE IMPLEMENTATION,
//                INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR
//                REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE
//                FROM CLAIMS OF INFRINGEMENT, IMPLIED WARRANTIES
//                OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
//                PURPOSE.
//
//                (c) Copyright 2008 Xilinx, Inc.
//                All rights reserved.
//

//
//  FRAME CHECK
//
//
//
//  Description: This module is a  pattern checker to test the Aurora
//               designs in hardware. The frames generated by FRAME_GEN
//               pass through the Aurora channel and arrive at the frame checker 
//               through the RX User interface. Every time an error is found in
//               the data recieved, the error count is incremented until it 
//               reaches its max value.

`timescale 1 ns / 10 ps
`define DLY #1


module aurora_RX_engine
(
    // User Interface
    RX_D,  
    RX_REM,     
    RX_SOF_N,       
    RX_EOF_N,
    RX_SRC_RDY_N,  

    // System Interface
    USER_CLK,       
    RESET,
    ERROR_COUNT,
	 
	 RX_DATA_VALID,
    RX_CLK_EN,
    RX_CLOCK,
    RX_DATA
  
);

//***********************************Port Declarations*******************************

   // User Interface
    input   [0:31]     RX_D;
    input   [0:1]      RX_REM;
    input              RX_SOF_N;
    input              RX_EOF_N;
    input              RX_SRC_RDY_N;
    
      // System Interface
    input              USER_CLK;
    input              RESET; 
    output  [0:7]      ERROR_COUNT;
	 
	 output RX_DATA_VALID;
    input RX_CLK_EN;
    input RX_CLOCK;
    output [31:0] RX_DATA;


//***************************Internal Register Declarations*************************** 

    reg                in_frame_r;
    //0:31]     data_r;
    reg                data_valid_r;
    //reg                error_detected_r;
    //reg     [0:8]      error_count_r;
    
 
//*********************************Wire Declarations**********************************
   
    wire               data_valid_c;
    wire               in_frame_c;
    wire               rem_valid_c;
    
    //wire               error_detected_c;


//*********************************Main Body of Code**********************************

wire empty;
assign RX_DATA_VALID = ~empty; 

aurora_FIFO RX (
.dout(RX_DATA),
.rd_clk(RX_CLOCK),
.rd_en(RX_CLK_EN),
.empty(empty),
.rst(RESET),
.wr_clk(USER_CLK),
.wr_en(data_valid_c),
.din(RX_D),
.full()
);
    


    //______________________________ Capture incoming data ___________________________    
    //Data is valid when RX_SRC_RDY_N is asserted and data is arriving within a frame
    assign  data_valid_c    =   in_frame_c && rem_valid_c && !RX_SRC_RDY_N;


    //Data is in a frame if it is a single cycle frame or a multi_cycle frame has started
    assign  in_frame_c  =   in_frame_r  ||  (!RX_SRC_RDY_N && !RX_SOF_N);
    
    
    //Start a multicycle frame when a frame starts without ending on the same cycle. End 
    //the frame when an EOF is detected
    always @(posedge USER_CLK)
        if(RESET)   
            in_frame_r  <=  `DLY    1'b0;
        else if(!in_frame_r && !RX_SOF_N && !RX_SRC_RDY_N && RX_EOF_N)
            in_frame_r  <=  `DLY    1'b1;
        else if(in_frame_r && !RX_SRC_RDY_N && !RX_EOF_N)
            in_frame_r  <=  `DLY    1'b0;
            
            
    //We expect rem to indicate a full word of data on the EOF cycle
    assign  rem_valid_c =   RX_EOF_N || (RX_REM == 2'd3);
                


    //Capture valid incoming data, right shifted 1 bit for comparison with the next valid
    //incoming data
  /*  always @(posedge USER_CLK)
        if(data_valid_c)    
            data_r  <=  `DLY    {RX_D[31],RX_D[0:30]};



    //Data in the data register is valid only if it was valid when captured and had no error
    always @(posedge USER_CLK)
        if(RESET)   data_valid_r    <=  `DLY    1'b0;
        else        data_valid_r    <=  `DLY    data_valid_c && !error_detected_c;



    
    //___________________________ Check incoming data for errors __________________________
         
    
    //An error is detected when valid data from the data register, when right shifted, does not match valid data
    //from the Aurora RX port
    assign  error_detected_c    =   data_valid_c && data_valid_r && (RX_D != data_r);   
    
    
    //We register the error_detected signal for use with the error counter logic
    always @(posedge USER_CLK)
        if(RESET)  
            error_detected_r    <=  `DLY    1'b0;
        else
            error_detected_r    <=  `DLY    error_detected_c;  

    
    
    //We count the total number of errors we detect. By keeping a count we make it less likely that we will miss
    //errors we did not directly observe. This counter must be reset when it reaches its max value
    always @(posedge USER_CLK)
        if(RESET)
            error_count_r       <=  `DLY    9'd0;
        else if(error_detected_r && !error_count_r[0] )
            error_count_r       <=  `DLY    error_count_r + 1;
            
    
    
    //Here we connect the lower 8 bits of the count (the MSbit is used only to check when the counter reaches
    //max value) to the module output
    assign  ERROR_COUNT =   error_count_r[1:8];*/
	 assign  ERROR_COUNT =   0;
    
    
endmodule           
